//=====================================================================
// Description:
// This header file
// Designer : extraordinary.h@sjtu.edu.cn
// Revision History
// V0 date:2024/12/14 Initial version, extraordinary.h@sjtu.edu.cn
//=====================================================================

//`define CHECK         // Enable the Assertion
`define DES           // Change the CODEC from XOR to DES
